--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   08:35:10 04/30/2020
-- Design Name:   
-- Module Name:   /home/ise/ael/registerbench_test.vhd
-- Project Name:  ael
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: registerbench
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY registerbench_test IS
END registerbench_test;
 
ARCHITECTURE behavior OF registerbench_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT registerbench
    PORT(
         ADDRA : IN  std_logic_vector(3 downto 0);
         ADDRB : IN  std_logic_vector(3 downto 0);
         ADDRW : IN  std_logic_vector(3 downto 0);
         W : IN  std_logic;
         DATA : IN  std_logic_vector(7 downto 0);
         RST : IN  std_logic;
         CLK : IN  std_logic;
         QA : OUT  std_logic_vector(7 downto 0);
         QB : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal ADDRA : std_logic_vector(3 downto 0) := (others => '0');
   signal ADDRB : std_logic_vector(3 downto 0) := (others => '0');
   signal ADDRW : std_logic_vector(3 downto 0) := (others => '0');
   signal W : std_logic := '0';
   signal DATA : std_logic_vector(7 downto 0) := (others => '0');
   signal RST : std_logic := '1';
   signal CLK : std_logic := '0';

 	--Outputs
   signal QA : std_logic_vector(7 downto 0);
   signal QB : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: registerbench PORT MAP (
          ADDRA => ADDRA,
          ADDRB => ADDRB,
          ADDRW => ADDRW,
          W => W,
          DATA => DATA,
          RST => RST,
          CLK => CLK,
          QA => QA,
          QB => QB
        );

   -- Clock process definitions
   CLK_process :process
   begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		ADDRW <= X"A" ; 
		W <= '1' ; 
		DATA <= X"64" ; 
		wait for 100 ns ; 
		ADDRA <= X"A" ;
		

      -- insert stimulus here 

      wait;
   end process;

END;
